* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
X0 a_891_413# a_193_47# a_975_413# VPB sky130_fd_pr__pfet_01v8  w= 0.42 l= 0.15
X1 a_1059_315# a_891_413# VGND VNB sky130_fd_pr__nfet_01v8      w= 0.65 l= 0.15
X2 a_466_413# a_27_47# a_561_413# VPB sky130_fd_pr__pfet_01v8   w= 0.42 l= 0.15
X3 a_634_159# a_27_47# a_891_413# VPB sky130_fd_pr__pfet_01v8   w= 0.42 l= 0.15
X4 a_381_47# a_193_47# a_466_413# VPB sky130_fd_pr__pfet_01v8   w= 0.42 l= 0.15
X5 VPWR D a_381_47# VPB sky130_fd_pr__pfet_01v8                 w= 0.42 l= 0.15
X6 VPWR a_466_413# a_634_159# VPB sky130_fd_pr__pfet_01v8       w= 0.75 l= 0.15
X7 VGND a_466_413# a_634_159# VNB sky130_fd_pr__nfet_01v8       w= 0.64 l= 0.15
X8 a_1017_47# a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8      w= 0.42 l= 0.15
X9 a_1059_315# a_891_413# VPWR VPB sky130_fd_pr__pfet_01v8      w= 1    l= 0.15
X10 a_561_413# a_634_159# VPWR VPB sky130_fd_pr__pfet_01v8      w= 0.42 l= 0.15
X11 VPWR a_1059_315# Q VPB sky130_fd_pr__pfet_01v8              w= 1    l= 0.15
X12 a_891_413# a_27_47# a_1017_47# VNB sky130_fd_pr__nfet_01v8  w= 0.36 l= 0.15
X13 a_634_159# a_193_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 w= 0.36 l= 0.15
X14 a_592_47# a_634_159# VGND VNB sky130_fd_pr__nfet_01v8       w= 0.42 l= 0.15
X15 a_466_413# a_193_47# a_592_47# VNB sky130_fd_pr__nfet_01v8  w= 0.36 l= 0.15
X16 VGND a_27_47# a_193_47# VNB sky130_fd_pr__nfet_01v8         w= 0.42 l= 0.15
X17 a_381_47# a_27_47# a_466_413# VNB sky130_fd_pr__nfet_01v8   w= 0.36 l= 0.15
X18 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8               w= 0.42 l= 0.15
X19 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8               w= 0.64 l= 0.15
X20 VPWR a_27_47# a_193_47# VPB sky130_fd_pr__pfet_01v8         w= 0.64 l= 0.15
X21 VGND D a_381_47# VNB sky130_fd_pr__nfet_01v8                w= 0.42 l= 0.15
X22 a_975_413# a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8     w= 0.42 l= 0.15
X23 VGND a_1059_315# Q VNB sky130_fd_pr__nfet_01v8              w= 0.65 l= 0.15
.ends