set ngbehavior=ltpsa

.lib "./libs/models/sky130.lib.spice" tt
.include "sky130_fd_sc_hd__dfxtp_1.spice"
.include "sky130_fd_sc_hd__inv_1.spice"

*.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
*.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q

xdfxtp0 clk d0 gnd gnd v2 v2 q0 sky130_fd_sc_hd__dfxtp_1
xdfxtp1 clk q0 gnd gnd v2 v2 q1 sky130_fd_sc_hd__dfxtp_1
xdfxtp2 clk q1 gnd gnd v2 v2 q2 sky130_fd_sc_hd__dfxtp_1
xdfxtp3 clk q2 gnd gnd v2 v2 q3 sky130_fd_sc_hd__dfxtp_1
xinv0 q3 gnd gnd v1 v1 out1 sky130_fd_sc_hd__inv_1

Vclk clk gnd pulse 0 1.8 0ns 0.1ns 0.1ns 1ns 2ns
Vin d0 gnd pulse 0 1.8 0.5ns 0.1ns 0.1ns 2ns 4ns
V1 v1 gnd dc 1.0V
V2 v2 gnd pulse 0 1.2 0.7ns 0.1ns 0.1ns 7ns 14ns
Vout out1 gnd

.tran 0.01n 24n
.control
run

plot V(clk)+12 V(d0)+10 V(q0)+8 V(q1)+6 V(q2)+4 V(q3)+2 V(out1)

*plot avg(-i(v1))*V(v1)
*plot avg(-i(v2))*V(v2)

.endc
.end

