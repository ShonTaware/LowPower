

.lib "./libs/models/sky130.lib.spice" tt
.include "sky130_fd_sc_hd__inv_1.spice"

xinv1 in1 gnd gnd v1 v1 o1 sky130_fd_sc_hd__inv_1
xinv2 o1 gnd gnd v2 v2 out1 sky130_fd_sc_hd__inv_1

V1 v1 gnd pulse 0.9 2.7 0ns 10ns 3ns 0ns 10ns
V2 v2 gnd dc 1.8V
Vout out1 gnd
*Vin in1 gnd pulse 0 1.8 0 0.1ns 0.1ns 2ns 4ns
Vin in1 gnd pulse 0 1.8 0.01ns 0.1ns 0.1ns 10ns 20ns

*.dc V2 0.5 1.5 0.1 V1 0.25 2.25 0.1 
*.dc V2 1.5 1.5 0.1 V1 0.75 2.25 0.1 
*.dc V1 0.9 2.7 0.1 

.tran 0.01n 20n
.control
run
plot V(v1)+10 V(v2)+8 V(in1)+6 V(o1)+3 V(out1)
plot avg(-i(v1))*V(v1)
plot avg(-i(v2))*V(v2)

*plot V(in1)+8 V(o1)+2 V(out1)
*plot V(v2)
*plot V(in1)
*plot V(out1)
*plot V(in1, out1)
.endc
.end

